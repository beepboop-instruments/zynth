----------------------------------------------------------------------------------
-- Company: beepboop
-- Engineer: Tyler Huddleston
-- 
-- Create Date: 03/22/2025
-- Design Name: Synthesizer Engine
-- Module Name: Synthesizer Package
-- Description: 
--   Contains constant and type definitions for the the synthesizer engine.
-- 
----------------------------------------------------------------------------------

library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;

package synth_pkg is
  constant SYNTH_ENG_REV  : std_logic_vector := x"00000003";
  constant SYNTH_ENG_DATE : std_logic_vector := x"04192025";

  -- memmory-mapped address definitions
  constant OFFSET_PULSE_WIDTH_REG  : std_logic_vector := "0000000"; --   0
  constant OFFSET_PULSE_REG        : std_logic_vector := "0000001"; --   1
  constant OFFSET_RAMP_REG         : std_logic_vector := "0000010"; --   2
  constant OFFSET_SAW_REG          : std_logic_vector := "0000011"; --   3
  constant OFFSET_TRI_REG          : std_logic_vector := "0000100"; --   4
  constant OFFSET_SINE_REG         : std_logic_vector := "0000101"; --   5
  constant OFFSET_GAIN_SHIFT_REG   : std_logic_vector := "0001000"; --  16
  constant OFFSET_GAIN_SCALE_REG   : std_logic_vector := "0001001"; --  17
  constant OFFSET_ADSR_ATTACK_AMT  : std_logic_vector := "0100000"; --  32
  constant OFFSET_ADSR_DECAY_AMT   : std_logic_vector := "0100001"; --  33
  constant OFFSET_ADSR_SUSTAIN_AMT : std_logic_vector := "0100010"; --  34
  constant OFFSET_ADSR_RELEASE_AMT : std_logic_vector := "0100011"; --  35
  constant OFFSET_COMP_ATTACK_AMT  : std_logic_vector := "0100100"; --  36
  constant OFFSET_COMP_RELEASE_AMT : std_logic_vector := "0100101"; --  37
  constant OFFSET_COMP_THRESHOLD   : std_logic_vector := "0100110"; --  38
  constant OFFSET_COMP_KNEE_WIDTH  : std_logic_vector := "0100111"; --  39
  constant OFFSET_COMP_KNEE_SLOPE  : std_logic_vector := "0101000"; --  40
  constant OFFSET_REV_REG          : std_logic_vector := "1111000"; -- 120
  constant OFFSET_DATE_REG         : std_logic_vector := "1111001"; -- 121
  constant OFFSET_WRAPBACK_REG     : std_logic_vector := "1111111"; -- 127

  -- vector size definitions
  constant WIDTH_WAVE_DATA   : natural := 16;
  constant WIDTH_PH_DATA     : natural := 32;
  constant WIDTH_NOTE_GAIN   : natural := 7;
  constant WIDTH_WAVE_GAIN   : natural := 7;
  constant WIDTH_OUT_DATA    : natural := 24;
  constant WIDTH_OUT_GAIN    : natural := 7;
  constant WIDTH_OUT_SHIFT   : natural := 5;
  constant WIDTH_PULSE_WIDTH : natural := 16;
  constant WIDTH_ADSR_COUNT  : natural := 20;
  constant WIDTH_ADSR_CC     : natural := 20;

  constant NUM_WFRMS       : natural := 5;
  constant NUM_NOTES       : natural := 128;
  constant I_LOWEST_NOTE   : natural := 0;
  constant I_HIGHEST_NOTE  : natural := I_LOWEST_NOTE + NUM_NOTES - 1;

  -- waveform indexes
  constant I_PULSE : natural := 0;
  constant I_RAMP  : natural := 1;
  constant I_SAW   : natural := 2;
  constant I_TRI   : natural := 3;
  constant I_SINE  : natural := 4;

  -- array data types
  type t_ph_inc_lut  is array (116 to 127) of unsigned(WIDTH_PH_DATA-1 downto 0);
  type t_ph_inc      is array (I_LOWEST_NOTE to I_HIGHEST_NOTE) of unsigned(WIDTH_PH_DATA-1 downto 0);
  type t_wave_data   is array (I_LOWEST_NOTE to I_HIGHEST_NOTE) of signed(WIDTH_WAVE_DATA-1 downto 0);
  type t_note_amp    is array (0 to 127) of unsigned(WIDTH_NOTE_GAIN-1 downto 0);
  type t_wfrm_amp    is array (0 to NUM_WFRMS-1) of unsigned(WIDTH_WAVE_GAIN-1 downto 0);
  type t_wfrm_ph     is array (0 to NUM_WFRMS-1) of unsigned(WIDTH_WAVE_DATA-1 downto 0);

  type t_adsr        is array (0 to 7) of unsigned(WIDTH_ADSR_COUNT-1 downto 0);
  type t_adsr_count  is array (I_LOWEST_NOTE to I_HIGHEST_NOTE) of unsigned(WIDTH_ADSR_COUNT-1 downto 0);
  type t_note_acc    is array (I_LOWEST_NOTE to I_HIGHEST_NOTE) of unsigned(WIDTH_ADSR_COUNT-1 downto 0);

end synth_pkg;

package body synth_pkg is
    -- No implementation needed for a package with only constants
end synth_pkg;
